library verilog;
use verilog.vl_types.all;
entity ALU_32bit_tb is
end ALU_32bit_tb;

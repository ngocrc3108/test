library verilog;
use verilog.vl_types.all;
entity RAM_tb is
end RAM_tb;

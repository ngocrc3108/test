library verilog;
use verilog.vl_types.all;
entity Processor_tb is
end Processor_tb;
